// sys.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module sys (
		input  wire        clk_clk,                            //                         clk.clk
		output wire        master_0_master_reset_reset,        //       master_0_master_reset.reset
		output wire [31:0] pin_out_external_connection_export, // pin_out_external_connection.export
		input  wire [31:0] pio_in_external_connection_export,  //  pio_in_external_connection.export
		input  wire        pulpino_0_config_testmode_i,        //            pulpino_0_config.testmode_i
		input  wire        pulpino_0_config_fetch_enable_i,    //                            .fetch_enable_i
		input  wire        pulpino_0_config_clock_gating_i,    //                            .clock_gating_i
		input  wire [31:0] pulpino_0_config_boot_addr_i,       //                            .boot_addr_i
		input  wire        reset_reset_n                       //                       reset.reset_n
	);

	wire  [31:0] pulpino_0_avalon_master_instr_readdata;                       // mm_interconnect_0:pulpino_0_avalon_master_instr_readdata -> pulpino_0:instr_rdata
	wire         pulpino_0_avalon_master_instr_waitrequest;                    // mm_interconnect_0:pulpino_0_avalon_master_instr_waitrequest -> pulpino_0:instr_busy
	wire  [31:0] pulpino_0_avalon_master_instr_address;                        // pulpino_0:instr_addr -> mm_interconnect_0:pulpino_0_avalon_master_instr_address
	wire         pulpino_0_avalon_master_instr_read;                           // pulpino_0:instr_read -> mm_interconnect_0:pulpino_0_avalon_master_instr_read
	wire         pulpino_0_avalon_master_instr_readdatavalid;                  // mm_interconnect_0:pulpino_0_avalon_master_instr_readdatavalid -> pulpino_0:instr_rvalid
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] pulpino_0_avalon_master_lsu_readdata;                         // mm_interconnect_1:pulpino_0_avalon_master_lsu_readdata -> pulpino_0:lsu_rdata
	wire         pulpino_0_avalon_master_lsu_waitrequest;                      // mm_interconnect_1:pulpino_0_avalon_master_lsu_waitrequest -> pulpino_0:lsu_busy
	wire  [31:0] pulpino_0_avalon_master_lsu_address;                          // pulpino_0:lsu_addr -> mm_interconnect_1:pulpino_0_avalon_master_lsu_address
	wire         pulpino_0_avalon_master_lsu_read;                             // pulpino_0:lsu_read -> mm_interconnect_1:pulpino_0_avalon_master_lsu_read
	wire   [3:0] pulpino_0_avalon_master_lsu_byteenable;                       // pulpino_0:lsu_be -> mm_interconnect_1:pulpino_0_avalon_master_lsu_byteenable
	wire         pulpino_0_avalon_master_lsu_readdatavalid;                    // mm_interconnect_1:pulpino_0_avalon_master_lsu_readdatavalid -> pulpino_0:lsu_rvalid
	wire   [1:0] pulpino_0_avalon_master_lsu_response;                         // mm_interconnect_1:pulpino_0_avalon_master_lsu_response -> pulpino_0:lsu_resp
	wire         pulpino_0_avalon_master_lsu_write;                            // pulpino_0:lsu_write -> mm_interconnect_1:pulpino_0_avalon_master_lsu_write
	wire  [31:0] pulpino_0_avalon_master_lsu_writedata;                        // pulpino_0:lsu_wdata -> mm_interconnect_1:pulpino_0_avalon_master_lsu_writedata
	wire         pulpino_0_avalon_master_lsu_writeresponsevalid;               // mm_interconnect_1:pulpino_0_avalon_master_lsu_writeresponsevalid -> pulpino_0:lsu_wrespvalid
	wire  [31:0] master_0_master_readdata;                                     // mm_interconnect_1:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                                  // mm_interconnect_1:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                      // master_0:master_address -> mm_interconnect_1:master_0_master_address
	wire         master_0_master_read;                                         // master_0:master_read -> mm_interconnect_1:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                   // master_0:master_byteenable -> mm_interconnect_1:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                                // mm_interconnect_1:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                        // master_0:master_write -> mm_interconnect_1:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                    // master_0:master_writedata -> mm_interconnect_1:master_0_master_writedata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_1_pin_out_s1_chipselect;                      // mm_interconnect_1:pin_out_s1_chipselect -> pin_out:chipselect
	wire  [31:0] mm_interconnect_1_pin_out_s1_readdata;                        // pin_out:readdata -> mm_interconnect_1:pin_out_s1_readdata
	wire   [1:0] mm_interconnect_1_pin_out_s1_address;                         // mm_interconnect_1:pin_out_s1_address -> pin_out:address
	wire         mm_interconnect_1_pin_out_s1_write;                           // mm_interconnect_1:pin_out_s1_write -> pin_out:write_n
	wire  [31:0] mm_interconnect_1_pin_out_s1_writedata;                       // mm_interconnect_1:pin_out_s1_writedata -> pin_out:writedata
	wire  [31:0] mm_interconnect_1_pio_in_s1_readdata;                         // pio_in:readdata -> mm_interconnect_1:pio_in_s1_readdata
	wire   [1:0] mm_interconnect_1_pio_in_s1_address;                          // mm_interconnect_1:pio_in_s1_address -> pio_in:address
	wire         mm_interconnect_1_onchip_memory2_0_s2_chipselect;             // mm_interconnect_1:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s2_readdata;               // onchip_memory2_0:readdata2 -> mm_interconnect_1:onchip_memory2_0_s2_readdata
	wire  [12:0] mm_interconnect_1_onchip_memory2_0_s2_address;                // mm_interconnect_1:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s2_byteenable;             // mm_interconnect_1:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	wire         mm_interconnect_1_onchip_memory2_0_s2_write;                  // mm_interconnect_1:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s2_writedata;              // mm_interconnect_1:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire         mm_interconnect_1_onchip_memory2_0_s2_clken;                  // mm_interconnect_1:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire  [31:0] mm_interconnect_1_pulpino_0_avalon_slave_debug_readdata;      // pulpino_0:debug_rdata -> mm_interconnect_1:pulpino_0_avalon_slave_debug_readdata
	wire         mm_interconnect_1_pulpino_0_avalon_slave_debug_waitrequest;   // pulpino_0:debug_busy -> mm_interconnect_1:pulpino_0_avalon_slave_debug_waitrequest
	wire  [14:0] mm_interconnect_1_pulpino_0_avalon_slave_debug_address;       // mm_interconnect_1:pulpino_0_avalon_slave_debug_address -> pulpino_0:debug_addr
	wire         mm_interconnect_1_pulpino_0_avalon_slave_debug_read;          // mm_interconnect_1:pulpino_0_avalon_slave_debug_read -> pulpino_0:debug_read
	wire         mm_interconnect_1_pulpino_0_avalon_slave_debug_readdatavalid; // pulpino_0:debug_rvalid -> mm_interconnect_1:pulpino_0_avalon_slave_debug_readdatavalid
	wire         mm_interconnect_1_pulpino_0_avalon_slave_debug_write;         // mm_interconnect_1:pulpino_0_avalon_slave_debug_write -> pulpino_0:debug_write
	wire  [31:0] mm_interconnect_1_pulpino_0_avalon_slave_debug_writedata;     // mm_interconnect_1:pulpino_0_avalon_slave_debug_writedata -> pulpino_0:debug_wdata
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] pulpino_0_interrupt_receiver_irq;                             // irq_mapper:sender_irq -> pulpino_0:irq_i
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:pulpino_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pulpino_0_reset_sink_reset_bridge_in_reset_reset, onchip_memory2_0:reset, pin_out:reset_n, pio_in:reset_n, pulpino_0:rst_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	altera_avalon_jtag_uart #(
		.readBufferDepth            (64),
		.readIRQThreshold           (8),
		.useRegistersForReadBuffer  (1),
		.useRegistersForWriteBuffer (1),
		.writeBufferDepth           (64),
		.writeIRQThreshold          (8),
		.printingMethod             (0),
		.FIFO_WIDTH                 (8),
		.WR_WIDTHU                  (6),
		.RD_WIDTHU                  (6),
		.write_le                   ("OFF"),
		.read_le                    ("OFF"),
		.HEX_WRITE_DEPTH_STR        (64),
		.HEX_READ_DEPTH_STR         (64),
		.legacySignalAllow          (0)
	) jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	sys_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   (master_0_master_reset_reset)    // master_reset.reset
	);

	sys_onchip_memory2_0 onchip_memory2_0 (
		.address     (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_1_onchip_memory2_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_1_onchip_memory2_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_1_onchip_memory2_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_1_onchip_memory2_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_1_onchip_memory2_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_1_onchip_memory2_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_1_onchip_memory2_0_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                                          //   clk1.clk
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	sys_pin_out pin_out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_pin_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pin_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pin_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pin_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pin_out_s1_readdata),   //                    .readdata
		.out_port   (pin_out_external_connection_export)       // external_connection.export
	);

	sys_pio_in pio_in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_1_pio_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_pio_in_s1_readdata), //                    .readdata
		.in_port  (pio_in_external_connection_export)     // external_connection.export
	);

	core_top #(
		.AXI_ADDR_WIDTH      (32),
		.AXI_DATA_WIDTH      (32),
		.AXI_ID_MASTER_WIDTH (10),
		.AXI_ID_SLAVE_WIDTH  (10),
		.AXI_USER_WIDTH      (0),
		.USE_ZERO_RISCY      (1),
		.RISCY_RV32F         (0),
		.ZERO_RV32M          (1),
		.ZERO_RV32E          (0)
	) pulpino_0 (
		.rst_n          (~rst_controller_reset_out_reset),                              //          reset_sink.reset_n
		.testmode_i     (pulpino_0_config_testmode_i),                                  //              config.testmode_i
		.fetch_enable_i (pulpino_0_config_fetch_enable_i),                              //                    .fetch_enable_i
		.clock_gating_i (pulpino_0_config_clock_gating_i),                              //                    .clock_gating_i
		.boot_addr_i    (pulpino_0_config_boot_addr_i),                                 //                    .boot_addr_i
		.clk            (clk_clk),                                                      //            clk_sink.clk
		.irq_i          (pulpino_0_interrupt_receiver_irq),                             //  interrupt_receiver.irq
		.instr_addr     (pulpino_0_avalon_master_instr_address),                        // avalon_master_instr.address
		.instr_rdata    (pulpino_0_avalon_master_instr_readdata),                       //                    .readdata
		.instr_read     (pulpino_0_avalon_master_instr_read),                           //                    .read
		.instr_rvalid   (pulpino_0_avalon_master_instr_readdatavalid),                  //                    .readdatavalid
		.instr_busy     (pulpino_0_avalon_master_instr_waitrequest),                    //                    .waitrequest
		.lsu_addr       (pulpino_0_avalon_master_lsu_address),                          //   avalon_master_lsu.address
		.lsu_rdata      (pulpino_0_avalon_master_lsu_readdata),                         //                    .readdata
		.lsu_read       (pulpino_0_avalon_master_lsu_read),                             //                    .read
		.lsu_rvalid     (pulpino_0_avalon_master_lsu_readdatavalid),                    //                    .readdatavalid
		.lsu_busy       (pulpino_0_avalon_master_lsu_waitrequest),                      //                    .waitrequest
		.lsu_write      (pulpino_0_avalon_master_lsu_write),                            //                    .write
		.lsu_be         (pulpino_0_avalon_master_lsu_byteenable),                       //                    .byteenable
		.lsu_wdata      (pulpino_0_avalon_master_lsu_writedata),                        //                    .writedata
		.lsu_resp       (pulpino_0_avalon_master_lsu_response),                         //                    .response
		.lsu_wrespvalid (pulpino_0_avalon_master_lsu_writeresponsevalid),               //                    .writeresponsevalid
		.debug_addr     (mm_interconnect_1_pulpino_0_avalon_slave_debug_address),       //  avalon_slave_debug.address
		.debug_rdata    (mm_interconnect_1_pulpino_0_avalon_slave_debug_readdata),      //                    .readdata
		.debug_read     (mm_interconnect_1_pulpino_0_avalon_slave_debug_read),          //                    .read
		.debug_rvalid   (mm_interconnect_1_pulpino_0_avalon_slave_debug_readdatavalid), //                    .readdatavalid
		.debug_busy     (mm_interconnect_1_pulpino_0_avalon_slave_debug_waitrequest),   //                    .waitrequest
		.debug_write    (mm_interconnect_1_pulpino_0_avalon_slave_debug_write),         //                    .write
		.debug_wdata    (mm_interconnect_1_pulpino_0_avalon_slave_debug_writedata)      //                    .writedata
	);

	sys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                          //                                  clk_0_clk.clk
		.pulpino_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // pulpino_0_reset_sink_reset_bridge_in_reset.reset
		.pulpino_0_avalon_master_instr_address            (pulpino_0_avalon_master_instr_address),            //              pulpino_0_avalon_master_instr.address
		.pulpino_0_avalon_master_instr_waitrequest        (pulpino_0_avalon_master_instr_waitrequest),        //                                           .waitrequest
		.pulpino_0_avalon_master_instr_read               (pulpino_0_avalon_master_instr_read),               //                                           .read
		.pulpino_0_avalon_master_instr_readdata           (pulpino_0_avalon_master_instr_readdata),           //                                           .readdata
		.pulpino_0_avalon_master_instr_readdatavalid      (pulpino_0_avalon_master_instr_readdatavalid),      //                                           .readdatavalid
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),    //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),      //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken)       //                                           .clken
	);

	sys_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.master_0_clk_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                               //   master_0_clk_reset_reset_bridge_in_reset.reset
		.pulpino_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // pulpino_0_reset_sink_reset_bridge_in_reset.reset
		.master_0_master_address                          (master_0_master_address),                                      //                            master_0_master.address
		.master_0_master_waitrequest                      (master_0_master_waitrequest),                                  //                                           .waitrequest
		.master_0_master_byteenable                       (master_0_master_byteenable),                                   //                                           .byteenable
		.master_0_master_read                             (master_0_master_read),                                         //                                           .read
		.master_0_master_readdata                         (master_0_master_readdata),                                     //                                           .readdata
		.master_0_master_readdatavalid                    (master_0_master_readdatavalid),                                //                                           .readdatavalid
		.master_0_master_write                            (master_0_master_write),                                        //                                           .write
		.master_0_master_writedata                        (master_0_master_writedata),                                    //                                           .writedata
		.pulpino_0_avalon_master_lsu_address              (pulpino_0_avalon_master_lsu_address),                          //                pulpino_0_avalon_master_lsu.address
		.pulpino_0_avalon_master_lsu_waitrequest          (pulpino_0_avalon_master_lsu_waitrequest),                      //                                           .waitrequest
		.pulpino_0_avalon_master_lsu_byteenable           (pulpino_0_avalon_master_lsu_byteenable),                       //                                           .byteenable
		.pulpino_0_avalon_master_lsu_read                 (pulpino_0_avalon_master_lsu_read),                             //                                           .read
		.pulpino_0_avalon_master_lsu_readdata             (pulpino_0_avalon_master_lsu_readdata),                         //                                           .readdata
		.pulpino_0_avalon_master_lsu_readdatavalid        (pulpino_0_avalon_master_lsu_readdatavalid),                    //                                           .readdatavalid
		.pulpino_0_avalon_master_lsu_write                (pulpino_0_avalon_master_lsu_write),                            //                                           .write
		.pulpino_0_avalon_master_lsu_writedata            (pulpino_0_avalon_master_lsu_writedata),                        //                                           .writedata
		.pulpino_0_avalon_master_lsu_response             (pulpino_0_avalon_master_lsu_response),                         //                                           .response
		.pulpino_0_avalon_master_lsu_writeresponsevalid   (pulpino_0_avalon_master_lsu_writeresponsevalid),               //                                           .writeresponsevalid
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.onchip_memory2_0_s2_address                      (mm_interconnect_1_onchip_memory2_0_s2_address),                //                        onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                        (mm_interconnect_1_onchip_memory2_0_s2_write),                  //                                           .write
		.onchip_memory2_0_s2_readdata                     (mm_interconnect_1_onchip_memory2_0_s2_readdata),               //                                           .readdata
		.onchip_memory2_0_s2_writedata                    (mm_interconnect_1_onchip_memory2_0_s2_writedata),              //                                           .writedata
		.onchip_memory2_0_s2_byteenable                   (mm_interconnect_1_onchip_memory2_0_s2_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s2_chipselect                   (mm_interconnect_1_onchip_memory2_0_s2_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s2_clken                        (mm_interconnect_1_onchip_memory2_0_s2_clken),                  //                                           .clken
		.pin_out_s1_address                               (mm_interconnect_1_pin_out_s1_address),                         //                                 pin_out_s1.address
		.pin_out_s1_write                                 (mm_interconnect_1_pin_out_s1_write),                           //                                           .write
		.pin_out_s1_readdata                              (mm_interconnect_1_pin_out_s1_readdata),                        //                                           .readdata
		.pin_out_s1_writedata                             (mm_interconnect_1_pin_out_s1_writedata),                       //                                           .writedata
		.pin_out_s1_chipselect                            (mm_interconnect_1_pin_out_s1_chipselect),                      //                                           .chipselect
		.pio_in_s1_address                                (mm_interconnect_1_pio_in_s1_address),                          //                                  pio_in_s1.address
		.pio_in_s1_readdata                               (mm_interconnect_1_pio_in_s1_readdata),                         //                                           .readdata
		.pulpino_0_avalon_slave_debug_address             (mm_interconnect_1_pulpino_0_avalon_slave_debug_address),       //               pulpino_0_avalon_slave_debug.address
		.pulpino_0_avalon_slave_debug_write               (mm_interconnect_1_pulpino_0_avalon_slave_debug_write),         //                                           .write
		.pulpino_0_avalon_slave_debug_read                (mm_interconnect_1_pulpino_0_avalon_slave_debug_read),          //                                           .read
		.pulpino_0_avalon_slave_debug_readdata            (mm_interconnect_1_pulpino_0_avalon_slave_debug_readdata),      //                                           .readdata
		.pulpino_0_avalon_slave_debug_writedata           (mm_interconnect_1_pulpino_0_avalon_slave_debug_writedata),     //                                           .writedata
		.pulpino_0_avalon_slave_debug_readdatavalid       (mm_interconnect_1_pulpino_0_avalon_slave_debug_readdatavalid), //                                           .readdatavalid
		.pulpino_0_avalon_slave_debug_waitrequest         (mm_interconnect_1_pulpino_0_avalon_slave_debug_waitrequest)    //                                           .waitrequest
	);

	sys_irq_mapper irq_mapper (
		.clk           (clk_clk),                          //       clk.clk
		.reset         (rst_controller_reset_out_reset),   // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),         // receiver0.irq
		.sender_irq    (pulpino_0_interrupt_receiver_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
